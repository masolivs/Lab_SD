-- biblioteca
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- entidade
entity maquinarefri is
    port (
        clk    : in  std_logic;
        moeda  : in  std_logic_vector(1 downto 0);
        r, c25, c50 : out std_logic
    );
end maquinarefri;
-- arquitetura
architecture rtl of maquinarefri is
    type state is (idle, e25c, e50c, e75c, e1, e125, d25c, d50c, d75c);
    signal currentstate, nextstate : state;
begin
    -- processo sincrono
    sync_proc: process(clk)
    begin
        if rising_edge(clk) then
            currentstate <= nextstate;
        end if;
    end process;
    -- processo combinacional
    comb_proc: process (currentstate, moeda)
    begin
        case currentstate is
            when idle =>
                r <= '0';
                c25 <= '0';
                c50 <= '0';
                if (moeda = "01") then
                    nextstate <= e25c;
                elsif (moeda = "10") then
                    nextstate <= e50c;
                else
                    nextstate <= idle;
                end if;
            when e25c =>
                r <= '0';
                c25 <= '0';
                c50 <= '0';
                if (moeda = "01") then
                    nextstate <= e50c;
                elsif (moeda = "10") then
                    nextstate <= e75c;
                elsif (moeda = "11") then
                    nextstate <= d25c;
                else
                    nextstate <= e25c;
                end if;
            when e50c =>
                r <= '0';
                c25 <= '0';
                c50 <= '0';
                if (moeda = "01") then
                    nextstate <= e75c;
                elsif (moeda = "10") then
                    nextstate <= e1;
                elsif (moeda = "11") then
                    nextstate <= d50c;
                else
                    nextstate <= e50c;
                end if;
            when e75c =>
                r <= '0';
                c25 <= '0';
                c50 <= '0';
                if (moeda = "01") then
                    nextstate <= e1;
                elsif (moeda = "10") then
                    nextstate <= e125;
                elsif (moeda = "11") then
                    nextstate <= d75c;
                else
                    nextstate <= e75c;
                end if;
            when e1 =>
                r <= '1';
                c25 <= '0';
                c50 <= '0';
                if (moeda = "01") then
                    nextstate <= e125;
                elsif (moeda = "10") then
                    nextstate <= e50c;
                else
                    nextstate <= idle;
                end if;
            when e125 =>
                r <= '1';
                c25 <= '1';
                c50 <= '0';
                if (moeda = "01") then
                    nextstate <= e25c;
                elsif (moeda = "10") then
                    nextstate <= e50c;
                else
                    nextstate <= idle;
                end if;
            when d25c =>
                r <= '0';
                c25 <= '1';
                c50 <= '0';
                if (moeda = "01") then
                    nextstate <= e25c;
                elsif (moeda = "10") then
                    nextstate <= e50c;
                else
                    nextstate <= idle;
                end if;
            when d50c =>
                r <= '0';
                c25 <= '0';
                c50 <= '1';
                if (moeda = "01") then
                    nextstate <= e25c;
                elsif (moeda = "10") then
                    nextstate <= e50c;
                else
                    nextstate <= idle;
                end if;
            when d75c =>
                r <= '0';
                c25 <= '1';
                c50 <= '1';
                if (moeda = "01") then
                    nextstate <= e25c;
                elsif (moeda = "10") then
                    nextstate <= e50c;
                else
                    nextstate <= idle;
                end if;
        end case;
    end process;
end rtl;
